`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oen,
    inout [`MPRJ_IO_PADS-8:0] analog_io,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    input   user_clock2    
);

core_top_wrapper 
core_wrapper ( 
    .vdda1(vdda1),	// User area 1 3.3V power
    .vdda2(vdda2),	// User area 2 3.3V power
    .vssa1(vssa1),	// User area 1 analog ground
    .vssa2(vssa2),	// User area 2 analog ground
    .vccd1(vccd1),	// User area 1 1.8V power
    .vccd2(vccd2),	// User area 2 1.8V power
    .vssd1(vssd1),	// User area 1 digital ground
    .vssd2(vssd2),	// User area 2 digital ground

    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),

        // MGMT SoC Wishbone Slave 
    .wbs_cyc_i  ( wbs_cyc_i     ),
    .wbs_stb_i  ( wbs_stb_i     ),
    .wbs_we_i   ( wbs_we_i      ),
    .wbs_sel_i  ( wbs_sel_i     ),
    .wbs_adr_i  ( wbs_adr_i     ),
    .wbs_dat_i  ( wbs_dat_i     ),
    .wbs_ack_o  ( wbs_ack_o     ),
    .wbs_dat_o  ( wbs_dat_o     ),

        // Logic Analyzer
    .la_data_in ( la_data_in    ),
    .la_data_out( la_data_out   ),
    .la_oen     ( la_oen        ),

        // IO Pads
    .io_in      ( io_in         ),
    .io_out     ( io_out        ),
    .io_oeb     ( io_oeb        ),
    .analog_io  ( analog_io     ),

    // Independent clock
    .user_clock2( mprj_clock2   )
);

endmodule	// user_project_wrapper
`default_nettype wire
