VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 597.600 2.670 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 597.600 157.690 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 597.600 172.870 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.230 597.600 188.510 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.870 597.600 204.150 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.510 597.600 219.790 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.690 597.600 234.970 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.330 597.600 250.610 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 597.600 266.250 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 597.600 281.890 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.790 597.600 297.070 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 597.600 17.850 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.430 597.600 312.710 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.070 597.600 328.350 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.250 597.600 343.530 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.890 597.600 359.170 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 597.600 374.810 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 597.600 390.450 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.350 597.600 405.630 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.990 597.600 421.270 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.630 597.600 436.910 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.270 597.600 452.550 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 597.600 33.490 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.450 597.600 467.730 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 483.090 597.600 483.370 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.730 597.600 499.010 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.910 597.600 514.190 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.550 597.600 529.830 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 545.190 597.600 545.470 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.830 597.600 561.110 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.010 597.600 576.290 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 597.600 49.130 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 597.600 64.310 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 597.600 79.950 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.310 597.600 95.590 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.950 597.600 111.230 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 597.600 126.410 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 597.600 142.050 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 597.600 7.730 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.470 597.600 162.750 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.110 597.600 178.390 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 597.600 193.570 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.930 597.600 209.210 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.570 597.600 224.850 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 597.600 240.490 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 255.390 597.600 255.670 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 271.030 597.600 271.310 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.670 597.600 286.950 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 302.310 597.600 302.590 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 597.600 22.910 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.490 597.600 317.770 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.130 597.600 333.410 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.770 597.600 349.050 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 363.950 597.600 364.230 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.590 597.600 379.870 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.230 597.600 395.510 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.870 597.600 411.150 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.050 597.600 426.330 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.690 597.600 441.970 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 597.600 457.610 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 597.600 38.550 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.510 597.600 472.790 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.150 597.600 488.430 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.790 597.600 504.070 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.430 597.600 519.710 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.610 597.600 534.890 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 550.250 597.600 550.530 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 565.890 597.600 566.170 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 581.530 597.600 581.810 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 597.600 54.190 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 597.600 69.830 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 597.600 85.010 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 597.600 100.650 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 597.600 116.290 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 597.600 131.930 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.830 597.600 147.110 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.510 597.600 12.790 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.530 597.600 167.810 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 597.600 183.450 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.810 597.600 199.090 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.990 597.600 214.270 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.630 597.600 229.910 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 245.270 597.600 245.550 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.910 597.600 261.190 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.090 597.600 276.370 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.730 597.600 292.010 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.370 597.600 307.650 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.150 597.600 28.430 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.550 597.600 322.830 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.190 597.600 338.470 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 353.830 597.600 354.110 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.470 597.600 369.750 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.650 597.600 384.930 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 400.290 597.600 400.570 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.930 597.600 416.210 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.570 597.600 431.850 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.750 597.600 447.030 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.390 597.600 462.670 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 597.600 43.610 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 478.030 597.600 478.310 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.210 597.600 493.490 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.850 597.600 509.130 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 524.490 597.600 524.770 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.130 597.600 540.410 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.310 597.600 555.590 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.950 597.600 571.230 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.590 597.600 586.870 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 597.600 59.250 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 597.600 74.890 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 597.600 90.530 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 597.600 105.710 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 597.600 121.350 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.710 597.600 136.990 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.350 597.600 152.630 600.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 2.400 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 2.400 300.520 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 597.600 74.840 600.000 75.440 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 591.650 597.600 591.930 600.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 597.600 224.440 600.000 225.040 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 596.710 597.600 596.990 600.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 597.600 374.720 600.000 375.320 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 2.400 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 597.600 524.320 600.000 524.920 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 2.400 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 594.320 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 594.320 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 7.565 594.320 587.605 ;
      LAYER met1 ;
        RECT 0.530 4.800 597.010 587.760 ;
      LAYER met2 ;
        RECT 0.560 597.320 2.110 597.600 ;
        RECT 2.950 597.320 7.170 597.600 ;
        RECT 8.010 597.320 12.230 597.600 ;
        RECT 13.070 597.320 17.290 597.600 ;
        RECT 18.130 597.320 22.350 597.600 ;
        RECT 23.190 597.320 27.870 597.600 ;
        RECT 28.710 597.320 32.930 597.600 ;
        RECT 33.770 597.320 37.990 597.600 ;
        RECT 38.830 597.320 43.050 597.600 ;
        RECT 43.890 597.320 48.570 597.600 ;
        RECT 49.410 597.320 53.630 597.600 ;
        RECT 54.470 597.320 58.690 597.600 ;
        RECT 59.530 597.320 63.750 597.600 ;
        RECT 64.590 597.320 69.270 597.600 ;
        RECT 70.110 597.320 74.330 597.600 ;
        RECT 75.170 597.320 79.390 597.600 ;
        RECT 80.230 597.320 84.450 597.600 ;
        RECT 85.290 597.320 89.970 597.600 ;
        RECT 90.810 597.320 95.030 597.600 ;
        RECT 95.870 597.320 100.090 597.600 ;
        RECT 100.930 597.320 105.150 597.600 ;
        RECT 105.990 597.320 110.670 597.600 ;
        RECT 111.510 597.320 115.730 597.600 ;
        RECT 116.570 597.320 120.790 597.600 ;
        RECT 121.630 597.320 125.850 597.600 ;
        RECT 126.690 597.320 131.370 597.600 ;
        RECT 132.210 597.320 136.430 597.600 ;
        RECT 137.270 597.320 141.490 597.600 ;
        RECT 142.330 597.320 146.550 597.600 ;
        RECT 147.390 597.320 152.070 597.600 ;
        RECT 152.910 597.320 157.130 597.600 ;
        RECT 157.970 597.320 162.190 597.600 ;
        RECT 163.030 597.320 167.250 597.600 ;
        RECT 168.090 597.320 172.310 597.600 ;
        RECT 173.150 597.320 177.830 597.600 ;
        RECT 178.670 597.320 182.890 597.600 ;
        RECT 183.730 597.320 187.950 597.600 ;
        RECT 188.790 597.320 193.010 597.600 ;
        RECT 193.850 597.320 198.530 597.600 ;
        RECT 199.370 597.320 203.590 597.600 ;
        RECT 204.430 597.320 208.650 597.600 ;
        RECT 209.490 597.320 213.710 597.600 ;
        RECT 214.550 597.320 219.230 597.600 ;
        RECT 220.070 597.320 224.290 597.600 ;
        RECT 225.130 597.320 229.350 597.600 ;
        RECT 230.190 597.320 234.410 597.600 ;
        RECT 235.250 597.320 239.930 597.600 ;
        RECT 240.770 597.320 244.990 597.600 ;
        RECT 245.830 597.320 250.050 597.600 ;
        RECT 250.890 597.320 255.110 597.600 ;
        RECT 255.950 597.320 260.630 597.600 ;
        RECT 261.470 597.320 265.690 597.600 ;
        RECT 266.530 597.320 270.750 597.600 ;
        RECT 271.590 597.320 275.810 597.600 ;
        RECT 276.650 597.320 281.330 597.600 ;
        RECT 282.170 597.320 286.390 597.600 ;
        RECT 287.230 597.320 291.450 597.600 ;
        RECT 292.290 597.320 296.510 597.600 ;
        RECT 297.350 597.320 302.030 597.600 ;
        RECT 302.870 597.320 307.090 597.600 ;
        RECT 307.930 597.320 312.150 597.600 ;
        RECT 312.990 597.320 317.210 597.600 ;
        RECT 318.050 597.320 322.270 597.600 ;
        RECT 323.110 597.320 327.790 597.600 ;
        RECT 328.630 597.320 332.850 597.600 ;
        RECT 333.690 597.320 337.910 597.600 ;
        RECT 338.750 597.320 342.970 597.600 ;
        RECT 343.810 597.320 348.490 597.600 ;
        RECT 349.330 597.320 353.550 597.600 ;
        RECT 354.390 597.320 358.610 597.600 ;
        RECT 359.450 597.320 363.670 597.600 ;
        RECT 364.510 597.320 369.190 597.600 ;
        RECT 370.030 597.320 374.250 597.600 ;
        RECT 375.090 597.320 379.310 597.600 ;
        RECT 380.150 597.320 384.370 597.600 ;
        RECT 385.210 597.320 389.890 597.600 ;
        RECT 390.730 597.320 394.950 597.600 ;
        RECT 395.790 597.320 400.010 597.600 ;
        RECT 400.850 597.320 405.070 597.600 ;
        RECT 405.910 597.320 410.590 597.600 ;
        RECT 411.430 597.320 415.650 597.600 ;
        RECT 416.490 597.320 420.710 597.600 ;
        RECT 421.550 597.320 425.770 597.600 ;
        RECT 426.610 597.320 431.290 597.600 ;
        RECT 432.130 597.320 436.350 597.600 ;
        RECT 437.190 597.320 441.410 597.600 ;
        RECT 442.250 597.320 446.470 597.600 ;
        RECT 447.310 597.320 451.990 597.600 ;
        RECT 452.830 597.320 457.050 597.600 ;
        RECT 457.890 597.320 462.110 597.600 ;
        RECT 462.950 597.320 467.170 597.600 ;
        RECT 468.010 597.320 472.230 597.600 ;
        RECT 473.070 597.320 477.750 597.600 ;
        RECT 478.590 597.320 482.810 597.600 ;
        RECT 483.650 597.320 487.870 597.600 ;
        RECT 488.710 597.320 492.930 597.600 ;
        RECT 493.770 597.320 498.450 597.600 ;
        RECT 499.290 597.320 503.510 597.600 ;
        RECT 504.350 597.320 508.570 597.600 ;
        RECT 509.410 597.320 513.630 597.600 ;
        RECT 514.470 597.320 519.150 597.600 ;
        RECT 519.990 597.320 524.210 597.600 ;
        RECT 525.050 597.320 529.270 597.600 ;
        RECT 530.110 597.320 534.330 597.600 ;
        RECT 535.170 597.320 539.850 597.600 ;
        RECT 540.690 597.320 544.910 597.600 ;
        RECT 545.750 597.320 549.970 597.600 ;
        RECT 550.810 597.320 555.030 597.600 ;
        RECT 555.870 597.320 560.550 597.600 ;
        RECT 561.390 597.320 565.610 597.600 ;
        RECT 566.450 597.320 570.670 597.600 ;
        RECT 571.510 597.320 575.730 597.600 ;
        RECT 576.570 597.320 581.250 597.600 ;
        RECT 582.090 597.320 586.310 597.600 ;
        RECT 587.150 597.320 591.370 597.600 ;
        RECT 592.210 597.320 596.430 597.600 ;
        RECT 0.560 2.680 596.980 597.320 ;
        RECT 1.110 2.400 1.190 2.680 ;
        RECT 2.030 2.400 2.570 2.680 ;
        RECT 3.410 2.400 3.490 2.680 ;
        RECT 4.330 2.400 4.870 2.680 ;
        RECT 5.710 2.400 6.250 2.680 ;
        RECT 7.090 2.400 7.170 2.680 ;
        RECT 8.010 2.400 8.550 2.680 ;
        RECT 9.390 2.400 9.930 2.680 ;
        RECT 10.770 2.400 10.850 2.680 ;
        RECT 11.690 2.400 12.230 2.680 ;
        RECT 13.070 2.400 13.610 2.680 ;
        RECT 14.450 2.400 14.530 2.680 ;
        RECT 15.370 2.400 15.910 2.680 ;
        RECT 16.750 2.400 17.290 2.680 ;
        RECT 18.130 2.400 18.210 2.680 ;
        RECT 19.050 2.400 19.590 2.680 ;
        RECT 20.430 2.400 20.970 2.680 ;
        RECT 21.810 2.400 21.890 2.680 ;
        RECT 22.730 2.400 23.270 2.680 ;
        RECT 24.110 2.400 24.650 2.680 ;
        RECT 25.490 2.400 25.570 2.680 ;
        RECT 26.410 2.400 26.950 2.680 ;
        RECT 27.790 2.400 28.330 2.680 ;
        RECT 29.170 2.400 29.250 2.680 ;
        RECT 30.090 2.400 30.630 2.680 ;
        RECT 31.470 2.400 32.010 2.680 ;
        RECT 32.850 2.400 32.930 2.680 ;
        RECT 33.770 2.400 34.310 2.680 ;
        RECT 35.150 2.400 35.690 2.680 ;
        RECT 36.530 2.400 36.610 2.680 ;
        RECT 37.450 2.400 37.990 2.680 ;
        RECT 38.830 2.400 38.910 2.680 ;
        RECT 39.750 2.400 40.290 2.680 ;
        RECT 41.130 2.400 41.670 2.680 ;
        RECT 42.510 2.400 42.590 2.680 ;
        RECT 43.430 2.400 43.970 2.680 ;
        RECT 44.810 2.400 45.350 2.680 ;
        RECT 46.190 2.400 46.270 2.680 ;
        RECT 47.110 2.400 47.650 2.680 ;
        RECT 48.490 2.400 49.030 2.680 ;
        RECT 49.870 2.400 49.950 2.680 ;
        RECT 50.790 2.400 51.330 2.680 ;
        RECT 52.170 2.400 52.710 2.680 ;
        RECT 53.550 2.400 53.630 2.680 ;
        RECT 54.470 2.400 55.010 2.680 ;
        RECT 55.850 2.400 56.390 2.680 ;
        RECT 57.230 2.400 57.310 2.680 ;
        RECT 58.150 2.400 58.690 2.680 ;
        RECT 59.530 2.400 60.070 2.680 ;
        RECT 60.910 2.400 60.990 2.680 ;
        RECT 61.830 2.400 62.370 2.680 ;
        RECT 63.210 2.400 63.750 2.680 ;
        RECT 64.590 2.400 64.670 2.680 ;
        RECT 65.510 2.400 66.050 2.680 ;
        RECT 66.890 2.400 67.430 2.680 ;
        RECT 68.270 2.400 68.350 2.680 ;
        RECT 69.190 2.400 69.730 2.680 ;
        RECT 70.570 2.400 71.110 2.680 ;
        RECT 71.950 2.400 72.030 2.680 ;
        RECT 72.870 2.400 73.410 2.680 ;
        RECT 74.250 2.400 74.790 2.680 ;
        RECT 75.630 2.400 75.710 2.680 ;
        RECT 76.550 2.400 77.090 2.680 ;
        RECT 77.930 2.400 78.010 2.680 ;
        RECT 78.850 2.400 79.390 2.680 ;
        RECT 80.230 2.400 80.770 2.680 ;
        RECT 81.610 2.400 81.690 2.680 ;
        RECT 82.530 2.400 83.070 2.680 ;
        RECT 83.910 2.400 84.450 2.680 ;
        RECT 85.290 2.400 85.370 2.680 ;
        RECT 86.210 2.400 86.750 2.680 ;
        RECT 87.590 2.400 88.130 2.680 ;
        RECT 88.970 2.400 89.050 2.680 ;
        RECT 89.890 2.400 90.430 2.680 ;
        RECT 91.270 2.400 91.810 2.680 ;
        RECT 92.650 2.400 92.730 2.680 ;
        RECT 93.570 2.400 94.110 2.680 ;
        RECT 94.950 2.400 95.490 2.680 ;
        RECT 96.330 2.400 96.410 2.680 ;
        RECT 97.250 2.400 97.790 2.680 ;
        RECT 98.630 2.400 99.170 2.680 ;
        RECT 100.010 2.400 100.090 2.680 ;
        RECT 100.930 2.400 101.470 2.680 ;
        RECT 102.310 2.400 102.850 2.680 ;
        RECT 103.690 2.400 103.770 2.680 ;
        RECT 104.610 2.400 105.150 2.680 ;
        RECT 105.990 2.400 106.530 2.680 ;
        RECT 107.370 2.400 107.450 2.680 ;
        RECT 108.290 2.400 108.830 2.680 ;
        RECT 109.670 2.400 110.210 2.680 ;
        RECT 111.050 2.400 111.130 2.680 ;
        RECT 111.970 2.400 112.510 2.680 ;
        RECT 113.350 2.400 113.430 2.680 ;
        RECT 114.270 2.400 114.810 2.680 ;
        RECT 115.650 2.400 116.190 2.680 ;
        RECT 117.030 2.400 117.110 2.680 ;
        RECT 117.950 2.400 118.490 2.680 ;
        RECT 119.330 2.400 119.870 2.680 ;
        RECT 120.710 2.400 120.790 2.680 ;
        RECT 121.630 2.400 122.170 2.680 ;
        RECT 123.010 2.400 123.550 2.680 ;
        RECT 124.390 2.400 124.470 2.680 ;
        RECT 125.310 2.400 125.850 2.680 ;
        RECT 126.690 2.400 127.230 2.680 ;
        RECT 128.070 2.400 128.150 2.680 ;
        RECT 128.990 2.400 129.530 2.680 ;
        RECT 130.370 2.400 130.910 2.680 ;
        RECT 131.750 2.400 131.830 2.680 ;
        RECT 132.670 2.400 133.210 2.680 ;
        RECT 134.050 2.400 134.590 2.680 ;
        RECT 135.430 2.400 135.510 2.680 ;
        RECT 136.350 2.400 136.890 2.680 ;
        RECT 137.730 2.400 138.270 2.680 ;
        RECT 139.110 2.400 139.190 2.680 ;
        RECT 140.030 2.400 140.570 2.680 ;
        RECT 141.410 2.400 141.950 2.680 ;
        RECT 142.790 2.400 142.870 2.680 ;
        RECT 143.710 2.400 144.250 2.680 ;
        RECT 145.090 2.400 145.630 2.680 ;
        RECT 146.470 2.400 146.550 2.680 ;
        RECT 147.390 2.400 147.930 2.680 ;
        RECT 148.770 2.400 149.310 2.680 ;
        RECT 150.150 2.400 150.230 2.680 ;
        RECT 151.070 2.400 151.610 2.680 ;
        RECT 152.450 2.400 152.530 2.680 ;
        RECT 153.370 2.400 153.910 2.680 ;
        RECT 154.750 2.400 155.290 2.680 ;
        RECT 156.130 2.400 156.210 2.680 ;
        RECT 157.050 2.400 157.590 2.680 ;
        RECT 158.430 2.400 158.970 2.680 ;
        RECT 159.810 2.400 159.890 2.680 ;
        RECT 160.730 2.400 161.270 2.680 ;
        RECT 162.110 2.400 162.650 2.680 ;
        RECT 163.490 2.400 163.570 2.680 ;
        RECT 164.410 2.400 164.950 2.680 ;
        RECT 165.790 2.400 166.330 2.680 ;
        RECT 167.170 2.400 167.250 2.680 ;
        RECT 168.090 2.400 168.630 2.680 ;
        RECT 169.470 2.400 170.010 2.680 ;
        RECT 170.850 2.400 170.930 2.680 ;
        RECT 171.770 2.400 172.310 2.680 ;
        RECT 173.150 2.400 173.690 2.680 ;
        RECT 174.530 2.400 174.610 2.680 ;
        RECT 175.450 2.400 175.990 2.680 ;
        RECT 176.830 2.400 177.370 2.680 ;
        RECT 178.210 2.400 178.290 2.680 ;
        RECT 179.130 2.400 179.670 2.680 ;
        RECT 180.510 2.400 181.050 2.680 ;
        RECT 181.890 2.400 181.970 2.680 ;
        RECT 182.810 2.400 183.350 2.680 ;
        RECT 184.190 2.400 184.730 2.680 ;
        RECT 185.570 2.400 185.650 2.680 ;
        RECT 186.490 2.400 187.030 2.680 ;
        RECT 187.870 2.400 187.950 2.680 ;
        RECT 188.790 2.400 189.330 2.680 ;
        RECT 190.170 2.400 190.710 2.680 ;
        RECT 191.550 2.400 191.630 2.680 ;
        RECT 192.470 2.400 193.010 2.680 ;
        RECT 193.850 2.400 194.390 2.680 ;
        RECT 195.230 2.400 195.310 2.680 ;
        RECT 196.150 2.400 196.690 2.680 ;
        RECT 197.530 2.400 198.070 2.680 ;
        RECT 198.910 2.400 198.990 2.680 ;
        RECT 199.830 2.400 200.370 2.680 ;
        RECT 201.210 2.400 201.750 2.680 ;
        RECT 202.590 2.400 202.670 2.680 ;
        RECT 203.510 2.400 204.050 2.680 ;
        RECT 204.890 2.400 205.430 2.680 ;
        RECT 206.270 2.400 206.350 2.680 ;
        RECT 207.190 2.400 207.730 2.680 ;
        RECT 208.570 2.400 209.110 2.680 ;
        RECT 209.950 2.400 210.030 2.680 ;
        RECT 210.870 2.400 211.410 2.680 ;
        RECT 212.250 2.400 212.790 2.680 ;
        RECT 213.630 2.400 213.710 2.680 ;
        RECT 214.550 2.400 215.090 2.680 ;
        RECT 215.930 2.400 216.470 2.680 ;
        RECT 217.310 2.400 217.390 2.680 ;
        RECT 218.230 2.400 218.770 2.680 ;
        RECT 219.610 2.400 220.150 2.680 ;
        RECT 220.990 2.400 221.070 2.680 ;
        RECT 221.910 2.400 222.450 2.680 ;
        RECT 223.290 2.400 223.830 2.680 ;
        RECT 224.670 2.400 224.750 2.680 ;
        RECT 225.590 2.400 226.130 2.680 ;
        RECT 226.970 2.400 227.050 2.680 ;
        RECT 227.890 2.400 228.430 2.680 ;
        RECT 229.270 2.400 229.810 2.680 ;
        RECT 230.650 2.400 230.730 2.680 ;
        RECT 231.570 2.400 232.110 2.680 ;
        RECT 232.950 2.400 233.490 2.680 ;
        RECT 234.330 2.400 234.410 2.680 ;
        RECT 235.250 2.400 235.790 2.680 ;
        RECT 236.630 2.400 237.170 2.680 ;
        RECT 238.010 2.400 238.090 2.680 ;
        RECT 238.930 2.400 239.470 2.680 ;
        RECT 240.310 2.400 240.850 2.680 ;
        RECT 241.690 2.400 241.770 2.680 ;
        RECT 242.610 2.400 243.150 2.680 ;
        RECT 243.990 2.400 244.530 2.680 ;
        RECT 245.370 2.400 245.450 2.680 ;
        RECT 246.290 2.400 246.830 2.680 ;
        RECT 247.670 2.400 248.210 2.680 ;
        RECT 249.050 2.400 249.130 2.680 ;
        RECT 249.970 2.400 250.510 2.680 ;
        RECT 251.350 2.400 251.890 2.680 ;
        RECT 252.730 2.400 252.810 2.680 ;
        RECT 253.650 2.400 254.190 2.680 ;
        RECT 255.030 2.400 255.570 2.680 ;
        RECT 256.410 2.400 256.490 2.680 ;
        RECT 257.330 2.400 257.870 2.680 ;
        RECT 258.710 2.400 259.250 2.680 ;
        RECT 260.090 2.400 260.170 2.680 ;
        RECT 261.010 2.400 261.550 2.680 ;
        RECT 262.390 2.400 262.470 2.680 ;
        RECT 263.310 2.400 263.850 2.680 ;
        RECT 264.690 2.400 265.230 2.680 ;
        RECT 266.070 2.400 266.150 2.680 ;
        RECT 266.990 2.400 267.530 2.680 ;
        RECT 268.370 2.400 268.910 2.680 ;
        RECT 269.750 2.400 269.830 2.680 ;
        RECT 270.670 2.400 271.210 2.680 ;
        RECT 272.050 2.400 272.590 2.680 ;
        RECT 273.430 2.400 273.510 2.680 ;
        RECT 274.350 2.400 274.890 2.680 ;
        RECT 275.730 2.400 276.270 2.680 ;
        RECT 277.110 2.400 277.190 2.680 ;
        RECT 278.030 2.400 278.570 2.680 ;
        RECT 279.410 2.400 279.950 2.680 ;
        RECT 280.790 2.400 280.870 2.680 ;
        RECT 281.710 2.400 282.250 2.680 ;
        RECT 283.090 2.400 283.630 2.680 ;
        RECT 284.470 2.400 284.550 2.680 ;
        RECT 285.390 2.400 285.930 2.680 ;
        RECT 286.770 2.400 287.310 2.680 ;
        RECT 288.150 2.400 288.230 2.680 ;
        RECT 289.070 2.400 289.610 2.680 ;
        RECT 290.450 2.400 290.990 2.680 ;
        RECT 291.830 2.400 291.910 2.680 ;
        RECT 292.750 2.400 293.290 2.680 ;
        RECT 294.130 2.400 294.670 2.680 ;
        RECT 295.510 2.400 295.590 2.680 ;
        RECT 296.430 2.400 296.970 2.680 ;
        RECT 297.810 2.400 298.350 2.680 ;
        RECT 299.190 2.400 299.270 2.680 ;
        RECT 300.110 2.400 300.650 2.680 ;
        RECT 301.490 2.400 301.570 2.680 ;
        RECT 302.410 2.400 302.950 2.680 ;
        RECT 303.790 2.400 304.330 2.680 ;
        RECT 305.170 2.400 305.250 2.680 ;
        RECT 306.090 2.400 306.630 2.680 ;
        RECT 307.470 2.400 308.010 2.680 ;
        RECT 308.850 2.400 308.930 2.680 ;
        RECT 309.770 2.400 310.310 2.680 ;
        RECT 311.150 2.400 311.690 2.680 ;
        RECT 312.530 2.400 312.610 2.680 ;
        RECT 313.450 2.400 313.990 2.680 ;
        RECT 314.830 2.400 315.370 2.680 ;
        RECT 316.210 2.400 316.290 2.680 ;
        RECT 317.130 2.400 317.670 2.680 ;
        RECT 318.510 2.400 319.050 2.680 ;
        RECT 319.890 2.400 319.970 2.680 ;
        RECT 320.810 2.400 321.350 2.680 ;
        RECT 322.190 2.400 322.730 2.680 ;
        RECT 323.570 2.400 323.650 2.680 ;
        RECT 324.490 2.400 325.030 2.680 ;
        RECT 325.870 2.400 326.410 2.680 ;
        RECT 327.250 2.400 327.330 2.680 ;
        RECT 328.170 2.400 328.710 2.680 ;
        RECT 329.550 2.400 330.090 2.680 ;
        RECT 330.930 2.400 331.010 2.680 ;
        RECT 331.850 2.400 332.390 2.680 ;
        RECT 333.230 2.400 333.770 2.680 ;
        RECT 334.610 2.400 334.690 2.680 ;
        RECT 335.530 2.400 336.070 2.680 ;
        RECT 336.910 2.400 337.450 2.680 ;
        RECT 338.290 2.400 338.370 2.680 ;
        RECT 339.210 2.400 339.750 2.680 ;
        RECT 340.590 2.400 340.670 2.680 ;
        RECT 341.510 2.400 342.050 2.680 ;
        RECT 342.890 2.400 343.430 2.680 ;
        RECT 344.270 2.400 344.350 2.680 ;
        RECT 345.190 2.400 345.730 2.680 ;
        RECT 346.570 2.400 347.110 2.680 ;
        RECT 347.950 2.400 348.030 2.680 ;
        RECT 348.870 2.400 349.410 2.680 ;
        RECT 350.250 2.400 350.790 2.680 ;
        RECT 351.630 2.400 351.710 2.680 ;
        RECT 352.550 2.400 353.090 2.680 ;
        RECT 353.930 2.400 354.470 2.680 ;
        RECT 355.310 2.400 355.390 2.680 ;
        RECT 356.230 2.400 356.770 2.680 ;
        RECT 357.610 2.400 358.150 2.680 ;
        RECT 358.990 2.400 359.070 2.680 ;
        RECT 359.910 2.400 360.450 2.680 ;
        RECT 361.290 2.400 361.830 2.680 ;
        RECT 362.670 2.400 362.750 2.680 ;
        RECT 363.590 2.400 364.130 2.680 ;
        RECT 364.970 2.400 365.510 2.680 ;
        RECT 366.350 2.400 366.430 2.680 ;
        RECT 367.270 2.400 367.810 2.680 ;
        RECT 368.650 2.400 369.190 2.680 ;
        RECT 370.030 2.400 370.110 2.680 ;
        RECT 370.950 2.400 371.490 2.680 ;
        RECT 372.330 2.400 372.870 2.680 ;
        RECT 373.710 2.400 373.790 2.680 ;
        RECT 374.630 2.400 375.170 2.680 ;
        RECT 376.010 2.400 376.090 2.680 ;
        RECT 376.930 2.400 377.470 2.680 ;
        RECT 378.310 2.400 378.850 2.680 ;
        RECT 379.690 2.400 379.770 2.680 ;
        RECT 380.610 2.400 381.150 2.680 ;
        RECT 381.990 2.400 382.530 2.680 ;
        RECT 383.370 2.400 383.450 2.680 ;
        RECT 384.290 2.400 384.830 2.680 ;
        RECT 385.670 2.400 386.210 2.680 ;
        RECT 387.050 2.400 387.130 2.680 ;
        RECT 387.970 2.400 388.510 2.680 ;
        RECT 389.350 2.400 389.890 2.680 ;
        RECT 390.730 2.400 390.810 2.680 ;
        RECT 391.650 2.400 392.190 2.680 ;
        RECT 393.030 2.400 393.570 2.680 ;
        RECT 394.410 2.400 394.490 2.680 ;
        RECT 395.330 2.400 395.870 2.680 ;
        RECT 396.710 2.400 397.250 2.680 ;
        RECT 398.090 2.400 398.170 2.680 ;
        RECT 399.010 2.400 399.550 2.680 ;
        RECT 400.390 2.400 400.930 2.680 ;
        RECT 401.770 2.400 401.850 2.680 ;
        RECT 402.690 2.400 403.230 2.680 ;
        RECT 404.070 2.400 404.610 2.680 ;
        RECT 405.450 2.400 405.530 2.680 ;
        RECT 406.370 2.400 406.910 2.680 ;
        RECT 407.750 2.400 408.290 2.680 ;
        RECT 409.130 2.400 409.210 2.680 ;
        RECT 410.050 2.400 410.590 2.680 ;
        RECT 411.430 2.400 411.970 2.680 ;
        RECT 412.810 2.400 412.890 2.680 ;
        RECT 413.730 2.400 414.270 2.680 ;
        RECT 415.110 2.400 415.190 2.680 ;
        RECT 416.030 2.400 416.570 2.680 ;
        RECT 417.410 2.400 417.950 2.680 ;
        RECT 418.790 2.400 418.870 2.680 ;
        RECT 419.710 2.400 420.250 2.680 ;
        RECT 421.090 2.400 421.630 2.680 ;
        RECT 422.470 2.400 422.550 2.680 ;
        RECT 423.390 2.400 423.930 2.680 ;
        RECT 424.770 2.400 425.310 2.680 ;
        RECT 426.150 2.400 426.230 2.680 ;
        RECT 427.070 2.400 427.610 2.680 ;
        RECT 428.450 2.400 428.990 2.680 ;
        RECT 429.830 2.400 429.910 2.680 ;
        RECT 430.750 2.400 431.290 2.680 ;
        RECT 432.130 2.400 432.670 2.680 ;
        RECT 433.510 2.400 433.590 2.680 ;
        RECT 434.430 2.400 434.970 2.680 ;
        RECT 435.810 2.400 436.350 2.680 ;
        RECT 437.190 2.400 437.270 2.680 ;
        RECT 438.110 2.400 438.650 2.680 ;
        RECT 439.490 2.400 440.030 2.680 ;
        RECT 440.870 2.400 440.950 2.680 ;
        RECT 441.790 2.400 442.330 2.680 ;
        RECT 443.170 2.400 443.710 2.680 ;
        RECT 444.550 2.400 444.630 2.680 ;
        RECT 445.470 2.400 446.010 2.680 ;
        RECT 446.850 2.400 447.390 2.680 ;
        RECT 448.230 2.400 448.310 2.680 ;
        RECT 449.150 2.400 449.690 2.680 ;
        RECT 450.530 2.400 450.610 2.680 ;
        RECT 451.450 2.400 451.990 2.680 ;
        RECT 452.830 2.400 453.370 2.680 ;
        RECT 454.210 2.400 454.290 2.680 ;
        RECT 455.130 2.400 455.670 2.680 ;
        RECT 456.510 2.400 457.050 2.680 ;
        RECT 457.890 2.400 457.970 2.680 ;
        RECT 458.810 2.400 459.350 2.680 ;
        RECT 460.190 2.400 460.730 2.680 ;
        RECT 461.570 2.400 461.650 2.680 ;
        RECT 462.490 2.400 463.030 2.680 ;
        RECT 463.870 2.400 464.410 2.680 ;
        RECT 465.250 2.400 465.330 2.680 ;
        RECT 466.170 2.400 466.710 2.680 ;
        RECT 467.550 2.400 468.090 2.680 ;
        RECT 468.930 2.400 469.010 2.680 ;
        RECT 469.850 2.400 470.390 2.680 ;
        RECT 471.230 2.400 471.770 2.680 ;
        RECT 472.610 2.400 472.690 2.680 ;
        RECT 473.530 2.400 474.070 2.680 ;
        RECT 474.910 2.400 475.450 2.680 ;
        RECT 476.290 2.400 476.370 2.680 ;
        RECT 477.210 2.400 477.750 2.680 ;
        RECT 478.590 2.400 479.130 2.680 ;
        RECT 479.970 2.400 480.050 2.680 ;
        RECT 480.890 2.400 481.430 2.680 ;
        RECT 482.270 2.400 482.810 2.680 ;
        RECT 483.650 2.400 483.730 2.680 ;
        RECT 484.570 2.400 485.110 2.680 ;
        RECT 485.950 2.400 486.490 2.680 ;
        RECT 487.330 2.400 487.410 2.680 ;
        RECT 488.250 2.400 488.790 2.680 ;
        RECT 489.630 2.400 489.710 2.680 ;
        RECT 490.550 2.400 491.090 2.680 ;
        RECT 491.930 2.400 492.470 2.680 ;
        RECT 493.310 2.400 493.390 2.680 ;
        RECT 494.230 2.400 494.770 2.680 ;
        RECT 495.610 2.400 496.150 2.680 ;
        RECT 496.990 2.400 497.070 2.680 ;
        RECT 497.910 2.400 498.450 2.680 ;
        RECT 499.290 2.400 499.830 2.680 ;
        RECT 500.670 2.400 500.750 2.680 ;
        RECT 501.590 2.400 502.130 2.680 ;
        RECT 502.970 2.400 503.510 2.680 ;
        RECT 504.350 2.400 504.430 2.680 ;
        RECT 505.270 2.400 505.810 2.680 ;
        RECT 506.650 2.400 507.190 2.680 ;
        RECT 508.030 2.400 508.110 2.680 ;
        RECT 508.950 2.400 509.490 2.680 ;
        RECT 510.330 2.400 510.870 2.680 ;
        RECT 511.710 2.400 511.790 2.680 ;
        RECT 512.630 2.400 513.170 2.680 ;
        RECT 514.010 2.400 514.550 2.680 ;
        RECT 515.390 2.400 515.470 2.680 ;
        RECT 516.310 2.400 516.850 2.680 ;
        RECT 517.690 2.400 518.230 2.680 ;
        RECT 519.070 2.400 519.150 2.680 ;
        RECT 519.990 2.400 520.530 2.680 ;
        RECT 521.370 2.400 521.910 2.680 ;
        RECT 522.750 2.400 522.830 2.680 ;
        RECT 523.670 2.400 524.210 2.680 ;
        RECT 525.050 2.400 525.130 2.680 ;
        RECT 525.970 2.400 526.510 2.680 ;
        RECT 527.350 2.400 527.890 2.680 ;
        RECT 528.730 2.400 528.810 2.680 ;
        RECT 529.650 2.400 530.190 2.680 ;
        RECT 531.030 2.400 531.570 2.680 ;
        RECT 532.410 2.400 532.490 2.680 ;
        RECT 533.330 2.400 533.870 2.680 ;
        RECT 534.710 2.400 535.250 2.680 ;
        RECT 536.090 2.400 536.170 2.680 ;
        RECT 537.010 2.400 537.550 2.680 ;
        RECT 538.390 2.400 538.930 2.680 ;
        RECT 539.770 2.400 539.850 2.680 ;
        RECT 540.690 2.400 541.230 2.680 ;
        RECT 542.070 2.400 542.610 2.680 ;
        RECT 543.450 2.400 543.530 2.680 ;
        RECT 544.370 2.400 544.910 2.680 ;
        RECT 545.750 2.400 546.290 2.680 ;
        RECT 547.130 2.400 547.210 2.680 ;
        RECT 548.050 2.400 548.590 2.680 ;
        RECT 549.430 2.400 549.970 2.680 ;
        RECT 550.810 2.400 550.890 2.680 ;
        RECT 551.730 2.400 552.270 2.680 ;
        RECT 553.110 2.400 553.650 2.680 ;
        RECT 554.490 2.400 554.570 2.680 ;
        RECT 555.410 2.400 555.950 2.680 ;
        RECT 556.790 2.400 557.330 2.680 ;
        RECT 558.170 2.400 558.250 2.680 ;
        RECT 559.090 2.400 559.630 2.680 ;
        RECT 560.470 2.400 561.010 2.680 ;
        RECT 561.850 2.400 561.930 2.680 ;
        RECT 562.770 2.400 563.310 2.680 ;
        RECT 564.150 2.400 564.230 2.680 ;
        RECT 565.070 2.400 565.610 2.680 ;
        RECT 566.450 2.400 566.990 2.680 ;
        RECT 567.830 2.400 567.910 2.680 ;
        RECT 568.750 2.400 569.290 2.680 ;
        RECT 570.130 2.400 570.670 2.680 ;
        RECT 571.510 2.400 571.590 2.680 ;
        RECT 572.430 2.400 572.970 2.680 ;
        RECT 573.810 2.400 574.350 2.680 ;
        RECT 575.190 2.400 575.270 2.680 ;
        RECT 576.110 2.400 576.650 2.680 ;
        RECT 577.490 2.400 578.030 2.680 ;
        RECT 578.870 2.400 578.950 2.680 ;
        RECT 579.790 2.400 580.330 2.680 ;
        RECT 581.170 2.400 581.710 2.680 ;
        RECT 582.550 2.400 582.630 2.680 ;
        RECT 583.470 2.400 584.010 2.680 ;
        RECT 584.850 2.400 585.390 2.680 ;
        RECT 586.230 2.400 586.310 2.680 ;
        RECT 587.150 2.400 587.690 2.680 ;
        RECT 588.530 2.400 589.070 2.680 ;
        RECT 589.910 2.400 589.990 2.680 ;
        RECT 590.830 2.400 591.370 2.680 ;
        RECT 592.210 2.400 592.750 2.680 ;
        RECT 593.590 2.400 593.670 2.680 ;
        RECT 594.510 2.400 595.050 2.680 ;
        RECT 595.890 2.400 596.430 2.680 ;
      LAYER met3 ;
        RECT 2.825 10.715 560.240 587.685 ;
      LAYER met4 ;
        RECT 21.040 10.640 560.240 587.760 ;
      LAYER met5 ;
        RECT 5.520 179.670 594.320 564.220 ;
  END
END user_proj_example
END LIBRARY

